`ifndef KEI_WATCHDOG_COV_SVH
`define KEI_WATCHDOG_COV_SVH

`include "kei_watchdog_cov.sv"


`endif //KEI_WATCHDOG_COV_SVH
