`ifndef KEI_WATCHDOG_CONFIG_SVH
`define KEI_WATCHDOG_CONFIG_SVH

`include "kei_watchdog_config.sv"

`endif
