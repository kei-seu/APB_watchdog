`ifndef KEI_WATCHDOG_TESTS_SVH
`define KEI_WATCHDOG_TESTS_SVH

`include "kei_watchdog_base_test.sv"
`include "kei_watchdog_apbacc_test.sv"
`include "kei_watchdog_regacc_test.sv"
`include "kei_watchdog_integration_test.sv"
`include "kei_watchdog_resen_test.sv"
`include "kei_watchdog_countdown_test.sv"
`include "kei_watchdog_disable_intr_test.sv"
`include "kei_watchdog_lock_test.sv"

`endif // KEI_WATCHDOG_TESTS_SVH
