`ifndef KEI_WATCHDOG_ELEMENT_SEQUENCES_LIB
`define KEI_WATCHDOG_ELEMENT_SEQUENCES_LIB

`include "kei_watchdog_base_element_sequence.sv"
`include "kei_watchdog_inrt_wait_clear.sv"
`include "kei_watchdog_loadcount.sv"
`include "kei_watchdog_reg_enable_inrt.sv"
`include "kei_watchdog_reg_enable_rst.sv"
`include "kei_watchdog_reg_disable_inrt.sv"
`include "kei_watchdog_reg_disable_rst.sv"



`endif  // KEI_WATCHDOG_ELEMENT_SEQUENCES_LIB
