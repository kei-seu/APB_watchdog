`ifndef KEI_WATCHDOG_REG
`define KEI_WATCHDOG_REG

`include "kei_watchdog_reg.sv"

`endif
