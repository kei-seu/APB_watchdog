`ifndef KEI_WATCHDOG_SEQ_LIB_SVH
`define KEI_WATCHDOG_SEQ_LIB_SVH

`include "kei_watchdog_element_sequences_lib.svh"
`include "kei_watchdog_base_virtual_sequence.sv"
`include "kei_watchdog_apbacc_virt_seq.sv"
`include "kei_watchdog_regacc_virt_seq.sv"
`include "kei_watchdog_integration_virt_seq.sv"
`include "kei_watchdog_resen_virt_seq.sv"
`include "kei_watchdog_countdown_virt_seq.sv"
`include "kei_watchdog_disable_intr_virt_seq.sv"

`endif 
